library ieee;

entity horas is
    port(
        ajuste          : in bit;
        modo            : in bit;
        minutos         : in bit;
        segundos        : in bit;
        hora            : out bit;
    )
    end horas;

    architecture hours of horas is
        begin
    
    end hours;