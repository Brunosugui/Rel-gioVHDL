library ieee;

entity minutos is
    port(
        segundos        : in bit;
        meio_segundos   : in bit;
        modo            : in bit;
        ajuste          : in bit;
        minuto          : out bit
    )
end minutos;

architecture minutes of minutos is
    begin
    
    end minutes;
